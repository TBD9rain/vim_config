//==============================================================================
//
//  Project         :   
//  File            :   
//  Version         :   v1.0
//  Title           :   
//                      
//  Description     :   
//                      
//  Addt'l info     :   
//  Version history :   
//
//  Author          :   
//  Email           :   
// 
//==============================================================================

module moduleName(
    //  IO PORT DECLARATIONS
    
);

//-----------------------
//  PARAMETER DEFINITIONS
//-----------------------



//---------------------
//  IO PORT DEFINITIONS
//---------------------



//----------------------
//  VARIABLE DEFINITIONS
//----------------------



//----------------
//  VERILOG CODING
//----------------



endmodule

