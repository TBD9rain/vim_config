//==============================================================================
//
//  Project         :   
//  File            :   
//  Version         :   v1.0
//  Title           :   
//                      
//  Description     :   
//                      
//  Addt'l info     :   
//  Version history :   
//
//  Author          :   
//  Email           :   
// 
//==============================================================================

module module_name(
    //  IO PORT DECLARATIONS
    
);

//-----------------------
//  PARAMETER DEFINITIONS
//-----------------------



//-----------------------
//  VARIABLES DEFINITIONS
//-----------------------



//----------------
//  VERILOG CODING
//----------------



endmodule
